interface mux_if ;
  logic [7:0] mux_in; 
  logic [2:0] mux_sel_in; 
  logic  mux_out; 
  

endinterface
